module not_gate(A, B);
    input wire A; 
    output wire B; 
    assign B = !A; 
endmodule

