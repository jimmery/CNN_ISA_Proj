// no simulations run. 
module max_decode(
    input clk, 
    input en, // turn on the max_decode.
    input [11:0] inst, 

    // how to do buffer stuff? 
)；

wire [3:0] in1_reg;
wire [3:0] in2_reg;
wire [3:0] dst_reg;

// represents the 32 max modules. 
reg [31:0] max_en;
reg [5:0] iterator;

assign in1_reg = inst[11:8];
assign in2_reg = inst[7:4];
assign dst_reg = inst[3:0];

reg [15:0] buffer [31:0] val;

reg [31:0] in1 [31:0] val1;
reg [31:0] in2 [31:0] val2;
wire [31:0] out [31:0] val3;

// define each module. 
max max_0(in1[0], in2[0], max_en[0], out[0]);
max max_1(in1[1], in2[1], max_en[1], out[1]);
max max_2(in1[2], in2[2], max_en[2], out[2]);
max max_3(in1[3], in2[3], max_en[3], out[3]);
max max_4(in1[4], in2[4], max_en[4], out[4]);
max max_5(in1[5], in2[5], max_en[5], out[5]);
max max_6(in1[6], in2[6], max_en[6], out[6]);
max max_7(in1[7], in2[7], max_en[7], out[7]);
max max_8(in1[8], in2[8], max_en[8], out[8]);
max max_9(in1[9], in2[9], max_en[9], out[9]);
max max_10(in1[10], in2[10], max_en[10], out[10]);
max max_11(in1[11], in2[11], max_en[11], out[11]);
max max_12(in1[12], in2[12], max_en[12], out[12]);
max max_13(in1[13], in2[13], max_en[13], out[13]);
max max_14(in1[14], in2[14], max_en[14], out[14]);
max max_15(in1[15], in2[15], max_en[15], out[15]);
max max_16(in1[16], in2[16], max_en[16], out[16]);
max max_17(in1[17], in2[17], max_en[17], out[17]);
max max_18(in1[18], in2[18], max_en[18], out[18]);
max max_19(in1[19], in2[19], max_en[19], out[19]);
max max_20(in1[20], in2[20], max_en[20], out[20]);
max max_21(in1[21], in2[21], max_en[21], out[21]);
max max_22(in1[22], in2[22], max_en[22], out[22]);
max max_23(in1[23], in2[23], max_en[23], out[23]);
max max_24(in1[24], in2[24], max_en[24], out[24]);
max max_25(in1[25], in2[25], max_en[25], out[25]);
max max_26(in1[26], in2[26], max_en[26], out[26]);
max max_27(in1[27], in2[27], max_en[27], out[27]);
max max_28(in1[28], in2[28], max_en[28], out[28]);
max max_29(in1[29], in2[29], max_en[29], out[29]);
max max_30(in1[30], in2[30], max_en[30], out[30]);
max max_31(in1[31], in2[31], max_en[31], out[31]);

initial
begin
  max_en = 32'b0;
  iterator = 5'b0;

  in1[0] = 32'b0;
  in1[1] = 32'b0;
  in1[2] = 32'b0;
  in1[3] = 32'b0;
  in1[4] = 32'b0;
  in1[5] = 32'b0;
  in1[6] = 32'b0;
  in1[7] = 32'b0;
  in1[8] = 32'b0;
  in1[9] = 32'b0;
  in1[10] = 32'b0;
  in1[11] = 32'b0;
  in1[12] = 32'b0;
  in1[13] = 32'b0;
  in1[14] = 32'b0;
  in1[15] = 32'b0;
  in1[16] = 32'b0;
  in1[17] = 32'b0;
  in1[18] = 32'b0;
  in1[19] = 32'b0;
  in1[20] = 32'b0;
  in1[21] = 32'b0;
  in1[22] = 32'b0;
  in1[23] = 32'b0;
  in1[24] = 32'b0;
  in1[25] = 32'b0;
  in1[26] = 32'b0;
  in1[27] = 32'b0;
  in1[28] = 32'b0;
  in1[29] = 32'b0;
  in1[30] = 32'b0;
  in1[31] = 32'b0;

  in2[0] = 32'b0;
  in2[1] = 32'b0;
  in2[2] = 32'b0;
  in2[3] = 32'b0;
  in2[4] = 32'b0;
  in2[5] = 32'b0;
  in2[6] = 32'b0;
  in2[7] = 32'b0;
  in2[8] = 32'b0;
  in2[9] = 32'b0;
  in2[10] = 32'b0;
  in2[11] = 32'b0;
  in2[12] = 32'b0;
  in2[13] = 32'b0;
  in2[14] = 32'b0;
  in2[15] = 32'b0;
  in2[16] = 32'b0;
  in2[17] = 32'b0;
  in2[18] = 32'b0;
  in2[19] = 32'b0;
  in2[20] = 32'b0;
  in2[21] = 32'b0;
  in2[22] = 32'b0;
  in2[23] = 32'b0;
  in2[24] = 32'b0;
  in2[25] = 32'b0;
  in2[26] = 32'b0;
  in2[27] = 32'b0;
  in2[28] = 32'b0;
  in2[29] = 32'b0;
  in2[30] = 32'b0;
  in2[31] = 32'b0;
end

always @(posedge clk)
begin
    iterator = 0; 
    max_en = 0;
    if (en) begin
        if (max_en[iterator])
            iterator = iterator + 1;
        end else begin
            in1[iterator] = buffer[in1_reg];
            in2[iterator] = buffer[in2_reg];
            max_en[iterator] = 1;

            buffer[dst_reg] = out[iterator];
            iterator = iterator + 1;
        end
    end
end
